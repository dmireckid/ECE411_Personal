import rv32i_types::*;

module mp2
(
    input clk,
    input rst,
    input pmem_resp,
    input [255:0] pmem_rdata,
    output logic pmem_read,
    output logic pmem_write,
    output rv32i_word pmem_address,
    output [255:0] pmem_wdata
);

logic [3:0] mem_byte_enable;
logic mem_read, mem_write, mem_resp;
rv32i_word mem_address, mem_wdata, mem_rdata;

// Keep cpu named `cpu` for RVFI Monitor
// Note: you have to rename your mp2 module to `cpu`
cpu cpu(.*);

// Keep cache named `cache` for RVFI Monitor
cache cache(.*);

// From MP0
//cacheline_adaptor cacheline_adaptor();

endmodule : mp2
